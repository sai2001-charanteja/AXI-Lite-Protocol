package axi_pkg;

	parameter ADDRESS_WIDTH = 16;
	parameter DATA_WIDTH    = 32;	
	parameter STRB_WIDTH    = 4;
	parameter DELAY_WIDTH    = 3;
	
	`include "axi_packet.sv"
endpackage
